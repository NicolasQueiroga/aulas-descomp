LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY decoderInstru IS
  PORT (
    opcode : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    saida : OUT STD_LOGIC_VECTOR(8 DOWNTO 0)
  );
END ENTITY;

ARCHITECTURE comportamento OF decoderInstru IS

  CONSTANT NOP : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0000";
  CONSTANT LDA : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0001";
  CONSTANT SOMA : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0010";
  CONSTANT SUB : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0011";
  CONSTANT LDI : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0100";
  CONSTANT STA : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0101";
  CONSTANT JMP : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0110";
  CONSTANT JEQ : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0110";
  CONSTANT CEQ : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0110";

BEGIN
  saida <= "0000XX000" WHEN opcode = NOP ELSE
    "000110010" WHEN opcode = LDA ELSE
    "000101010" WHEN opcode = SOMA ELSE
    "000100010" WHEN opcode = SUB ELSE
    "001110000" WHEN opcode = LDI ELSE
    "00X0XX001" WHEN opcode = STA ELSE
	 "10X0XX000" WHEN opcode = JMP ELSE
	 "01X0XX000" WHEN opcode = JEQ ELSE
	 "000000100" WHEN opcode = CEQ ELSE
    "000000000"; -- NOP para os opcodes Indefinidos
END ARCHITECTURE;